module calc(input wire clk,
            input wire btnac,
            input wire btnl,
            input wire btnr,
            input wire btnc,
            input wire btnd,
            input wire [15:0] sw,
            output wire [15:0] led);

    

endmodule
